module zpu_rom(
	input clk,
	input [addr_width-1:0] addr,
	output [7:0] dout);
	parameter addr_width = 8;
	reg [7:0] dout;
	reg [7:0] dout_rom0;
SB_ROM512x8 #(
.INIT_0(256'h80DA0B80C0A8808C0C0B0B0B0BA00881),
.INIT_1(256'h050B0B0B0BA00C0B0B0B0B8004000000),
.INIT_2(256'h00000001000000000000000000000000),
.INIT_3(256'h00000000000000900000000000000090),
.INIT_4(256'h0300D080C27F0000B012D080C27F0000),
.INIT_5(256'h2813D080C27F00001013D080C27F0300),
.INIT_6(256'h1005EF020100000065000D28FC0700C0),
.INIT_7(256'h5004EF0201000000700AD080C27F0000),
.INIT_8(256'h00FFEE0201000000700AD080C27F0000),
.INIT_9(256'h10FEEE0201000000D008D080C27F0000),
.INIT_A(256'h9009D080C27F00009405D080C27F0000),
.INIT_B(256'h5004EF0201000000A009D080C27F0000),
.INIT_C(256'h30FDEE02010000000006D080C27F0000),
.INIT_D(256'hE000EF0201000000F00AD080C27F0000),
.INIT_E(256'h2E006F757466696C653E2029207C2028),
.INIT_F(256'h1005EF02010000000000000000000090)
) _rom0 (
.RDATA(dout_rom0),
.RADDR(addr[8:0]),
.RCLK(clk), .RCLKE(1'b1), .RE(1'b1)
);
always @(posedge clk) begin
	dout <= dout_rom0;
end
endmodule
